`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:03:38 04/29/2014 
// Design Name: 
// Module Name:    Anti_jitter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Anti_jitter(input wire clk, 
						 input wire [3:0] button,
						 input wire [7:0] SW, 
						 output reg [3:0]button_out,
						 output reg [3:0]button_pulse,
						 output reg [7:0] SW_OK,
						 output reg rst

						);
	 
endmodule
